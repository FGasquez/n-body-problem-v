module main

import solver
import animation
import gx
import benchmark

struct BodiesContainer {
mut:
	bodies []solver.Body
	to_draw [][]solver.Body
}

fn main() {
	threads_count := 3
	mut threads := []thread{cap: threads_count}
	mut to_draw := [][]solver.Body{}
	requests := chan solver.BodyRequest{}
	results := chan solver.Body{}
	finished := chan bool{}

	delta := 0.001
	iterations_count := 500000
	g := 9.8

	mut bodies := [
		solver.Body{
			id: 0
			mass: 50.0
			color: gx.red
			unamovable: false
			pos: solver.Vector{
				x: 10.0
				y: 30.0
				z: 0.0
			}
			vel: solver.Vector{
				x: 0.0
				y: 0.0
				z: 0.0
			}
		},
		solver.Body{
			id: 1
			mass: 4.0
			color: gx.green
			unamovable: false
			pos: solver.Vector{
				x: 10.0
				y: 70.0
				z: 0.0
			}
			vel: solver.Vector{
				x: 3.5
				y: 0.0
				z: 0.0
			}
		},
		solver.Body{
			id: 2
			mass: 5.0
			color: gx.yellow
			unamovable: false
			pos: solver.Vector{
				x: -30.0
				y: -30.0
				z: 0.0
			}
			vel: solver.Vector{
				x: -2.0
				y: 2.0
				z: 0.0
			}
		},
		solver.Body{
			id: 3
			mass: 5.0
			color: gx.yellow
			unamovable: false
			pos: solver.Vector{
				x: -30.0
				y: -30.0
				z: 0.0
			}
			vel: solver.Vector{
				x: -2.0
				y: 2.0
				z: 0.0
			}
		},
			solver.Body{
			id: 4
			mass: 5.0
			color: gx.yellow
			unamovable: false
			pos: solver.Vector{
				x: -30.0
				y: -30.0
				z: 0.0
			}
			vel: solver.Vector{
				x: -2.0
				y: 2.0
				z: 0.0
			}
		},
			solver.Body{
			id: 5
			mass: 5.0
			color: gx.yellow
			unamovable: false
			pos: solver.Vector{
				x: -30.0
				y: -30.0
				z: 0.0
			}
			vel: solver.Vector{
				x: -2.0
				y: 2.0
				z: 0.0
			}
		}
	]

	to_draw << bodies.clone()

	mut container := &BodiesContainer{
		bodies: bodies
		to_draw: to_draw
	}

	mut bmark := benchmark.start()

	for i in 0 .. threads_count {
		threads << go solver.worker(requests, results, g, delta, i)
	}

	// go results_worker(mut container, results, finished)

	for _ in 0 .. iterations_count {
		println('x')
		prev_state := container.bodies.clone()
		for i in 0 .. container.bodies.len {
			requests <- solver.BodyRequest{
				body: prev_state[i]
				previous_state: prev_state
				id: i
			}
		}

		for i in 0 .. container.bodies.len {
			container.bodies[i] = <-results
		}
	}
	// for _ in 0 .. iterations_count {
	// 	prev_state := container.bodies.clone()
	// 	requests <- solver.BodyRequest{
	// 		body: prev_state[0]
	// 		previous_state: [prev_state[1], prev_state[2]]
	// 	}
	// 	requests <- solver.BodyRequest{
	// 		body: prev_state[1]
	// 		previous_state: [prev_state[0], prev_state[2]]
	// 	}
	// 	requests <- solver.BodyRequest{
	// 		body: prev_state[2]
	// 		previous_state: [prev_state[0], prev_state[1]]
	// 	}
	// 	_ := <- finished or { break }
	// }

	requests.close()
	threads.wait()

	finished.close()
	results.close()
	
	bmark.measure(@FN)

	animation.start(container.to_draw)
}

fn results_worker(mut container BodiesContainer, results chan solver.Body, finished chan bool) {
	mut i := 0
	for {
		res := <-results or { break }
		container.bodies[res.id] = res
		if i == container.bodies.len -1 {
			container.to_draw << container.bodies.clone()
			finished <- true
			i = -1
		}
		i++
	}
}
